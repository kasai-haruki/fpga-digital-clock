module CLOCK_ALL(CLK, RESET, LED, SA, btn_switch, btn_display, btn_inc); 
input CLK, RESET, btn_switch, btn_display, btn_inc; 
output [7:0] LED; 
output [3:0] SA; 
 
reg [26:0] tmp_count; 

wire [3:0] SEC_CNT10; 
wire [3:0] SEC_CNT6; 
wire [3:0] MIN_CNT10; 
wire [3:0] MIN_CNT6; 
wire [3:0] HOU_CNT10; 
wire [3:0] HOU_CNT3; 
wire [3:0] CNT_1, CNT_2, CNT_3, CNT_4, CNT; 
wire ENABLE, ENABLE_kHz; 
wire [7:0] L1, L2, L3, L4; 
wire CARRY, CARRY_2, CARRY_3, CARRY_4, CARRY_5, CARRY_6, is_leap, TOP_MODE, DIS_MODE, SET_MODE, INC_MODE;
wire [7:0] month;
wire [11:0] year;
//wire [15:0] WEEKDAY_LED;
wire [3:0] DAY_CNT10, DAY_CNT4, MON_CNT10, MON_CNT2, YEA_CNT10_1, YEA_CNT10_2, YEA_CNT2, week_day;
wire [4:0] TOP_CURRENT_STATE;
wire [6:0] DIS_CURRENT_STATE, SET_CURRENT_STATE;
assign month = {MON_CNT2, MON_CNT10};
assign year = {YEA_CNT2, YEA_CNT10_2, YEA_CNT10_1};

parameter SEC1_MAX = 125000000; // 125MHz 
 
CNT60 i0(.CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .CARRY_in(1'b1), .CARRY_out(CARRY), .INC_MODE(INC_MODE),
           .CNT10(SEC_CNT10), .CNT6(SEC_CNT6), .SET_CURRENT_STATE({SET_CURRENT_STATE[6], SET_CURRENT_STATE[0]})); 
DECODER7 i1(.COUNT(CNT), .LED(LED), .TOP_CURRENT_STATE(TOP_CURRENT_STATE[0]), .DIS_CURRENT_STATE(DIS_CURRENT_STATE[3:2]), .SA(SA)); 
CNT60 i2(.CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .CARRY_in(CARRY), .CARRY_out(CARRY_2),  .INC_MODE(INC_MODE),
           .CNT10(MIN_CNT10), .CNT6(MIN_CNT6), .SET_CURRENT_STATE({SET_CURRENT_STATE[5], SET_CURRENT_STATE[0]})); 
DCOUNT i3(.CLK(CLK), .ENABLE(ENABLE_kHz), .L1(CNT_1), .L2(CNT_2), 
          .L3(CNT_3), .L4(CNT_4), .SA(SA), .L(CNT)); 
CNT24 i4(.CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .CARRY_in(CARRY_2), .CARRY_out(CARRY_3), .INC_MODE(INC_MODE),
           .CNT10(HOU_CNT10), .CNT3(HOU_CNT3), .SET_CURRENT_STATE({SET_CURRENT_STATE[4], SET_CURRENT_STATE[0]}));  
SEC1 #(.SEC1_MAX(SEC1_MAX)) i5(.CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .ENABLE_kHz(ENABLE_kHz));
CNT_DAY i6(     .CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .CARRY_in(CARRY_3), .CARRY_out(CARRY_4), .INC_MODE(INC_MODE),
                .CNT10(DAY_CNT10), .CNT4(DAY_CNT4), .month(month), .is_leap(is_leap), .SET_CURRENT_STATE({SET_CURRENT_STATE[3], SET_CURRENT_STATE[0]})); 
CNT_MONTH i7(   .CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .CARRY_in(CARRY_4), .CARRY_out(CARRY_5), .INC_MODE(INC_MODE),
                .CNT10(MON_CNT10), .CNT2(MON_CNT2), .SET_CURRENT_STATE({SET_CURRENT_STATE[2], SET_CURRENT_STATE[0]}));  
CNT_YEAR i8(    .CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .CARRY_in(CARRY_5), .CARRY_out(CARRY_6), .INC_MODE(INC_MODE),
                .CNT10(YEA_CNT10_1), .CNT10_2(YEA_CNT10_2), .CNT2(YEA_CNT2), .SET_CURRENT_STATE({SET_CURRENT_STATE[1], SET_CURRENT_STATE[0]}));    
leap_year i9(   .year_bcd(year), .is_leap(is_leap));
//LED_WEEK i10(    .week_day(week_day), .LED(WEEKDAY_LED));
weekday_calc i10(.year_bcd(year), .month_bcd(month), .day_bcd({DAY_CNT4, DAY_CNT10}), .clk(CLK), .weekday(week_day));
MSE i11(.CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .MODE(TOP_MODE), .MODE_IN(btn_switch));
MAIN_MODE i12(.CLK(CLK), .RESET(RESET), .MODE(TOP_MODE), .CURRENT_STATE(TOP_CURRENT_STATE));
MSE i13(.CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .MODE(DIS_MODE), .MODE_IN(btn_display));
DIS_MODE i14(.CLK(CLK), .RESET(RESET), .MODE(DIS_MODE), .CURRENT_STATE(DIS_CURRENT_STATE), .main_state_active(TOP_CURRENT_STATE[0]));
MSE i15(.CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .MODE(SET_MODE), .MODE_IN(btn_display));
SET_MODE i16(.CLK(CLK), .RESET(RESET), .MODE(SET_MODE), .CURRENT_STATE(SET_CURRENT_STATE), .main_state_active(TOP_CURRENT_STATE[1]));
MSE i17(.CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .MODE(INC_MODE), .MODE_IN(btn_inc));
display_switch i18(     .TOP_CURRENT_STATE(TOP_CURRENT_STATE[1:0]), .DIS_CURRENT_STATE(DIS_CURRENT_STATE), .SET_CURRENT_STATE(SET_CURRENT_STATE),
                        .SEC_CNT10(SEC_CNT10), .SEC_CNT6(SEC_CNT6), .MIN_CNT10(MIN_CNT10), .MIN_CNT6(MIN_CNT6),
                        .HOU_CNT10(HOU_CNT10), .HOU_CNT3(HOU_CNT3), .DAY_CNT10(DAY_CNT10), .DAY_CNT4(DAY_CNT4), .week_day(week_day),
                        .MON_CNT10(MON_CNT10), .MON_CNT2(MON_CNT2), .YEA_CNT10_1(YEA_CNT10_1), .YEA_CNT10_2(YEA_CNT10_2), .YEA_CNT2(YEA_CNT2),
                        .C1_out(CNT_1), .C2_out(CNT_2), .C3_out(CNT_3), .C4_out(CNT_4));                
 
endmodule 